spice

*.options trace
v1 n1 0 pulse iv=0 pv=1 rise=1m delay=1 width=3 fall=1m
c1 n2 0 1
r1 n1 n2 1

.print tran v(nodes) method(c1) disc(nodes) hidden(0) event(v1)
.tran 0 2 2 trace=a

.stat

.options method traponly
.tran 0 2 2 trace=a

.stat
.end
