spice
v1 1 0 dc a ac b
.list
