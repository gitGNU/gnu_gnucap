spice

*.options trace
v1 n1 0 pulse iv=0 pv=1 rise=1m delay=1m width=3m fall=5m
c1 n2 0 200n
r1 n1 n2 1k

.print tran v(nodes) method(c1) disc(nodes) hidden(0) event(v1)
.tran 0 20m 20m trace=a

.stat

.options method traponly
.tran 0 20m 20m trace=a

.stat
.end
